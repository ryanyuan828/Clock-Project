LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_UNSIGNED.ALL;

ENTITY CALENDAR IS
PORT(
	CLK_100:IN STD_LOGIC;
	SETIN,CLRIN,RUNIN,ADDIN: IN STD_LOGIC;
	SET_NUM:IN STD_LOGIC_VECTOR(2 DOWNTO 0);
	MODE_NUM: IN STD_LOGIC_VECTOR(2 DOWNTO 0);
	
	CAL_E5,CAL_E4,CAL_E3,CAL_E2,CAL_E1,CAL_E0: INOUT STD_LOGIC_VECTOR(3 DOWNTO 0);
	CAL_D5,CAL_D4,CAL_D3,CAL_D2,CAL_D1,CAL_D0: INOUT STD_LOGIC_VECTOR(3 DOWNTO 0);
	CAL_START: OUT STD_LOGIC;
	CAL_ADD: IN STD_LOGIC
);
END ENTITY CALENDAR;

ARCHITECTURE BEHAVE OF CALENDAR IS
SIGNAL CAL_E5R,CAL_E4R,CAL_E3R,CAL_E2R,CAL_E1R,CAL_E0R: STD_LOGIC_VECTOR(3 DOWNTO 0);
SIGNAL CAL_D5R,CAL_D4R,CAL_D3R,CAL_D2R,CAL_D1R,CAL_D0R: STD_LOGIC_VECTOR(3 DOWNTO 0);
SIGNAL START: STD_LOGIC:='0';
SIGNAL CLR: STD_LOGIC:='1';
SIGNAL RUN,ADD: STD_LOGIC;

BEGIN
CAL_E5<=CAL_E5R;
CAL_E4<=CAL_E4R;
CAL_E3<=CAL_E3R;
CAL_E2<=CAL_E2R;
CAL_E1<=CAL_E1R;
CAL_E0<=CAL_E0R;

CAL_D5<=CAL_D5R;
CAL_D4<=CAL_D4R;
CAL_D3<=CAL_D3R;
CAL_D2<=CAL_D2R;
CAL_D1<=CAL_D1R;
CAL_D0<=CAL_D0R;
CAL_START<=START;

ADD1:PROCESS(ADDIN)
BEGIN
	IF(MODE_NUM="001" AND ADDIN='1') THEN
		ADD<='1';
	ELSE
		ADD<='0';
	END IF;
END PROCESS ADD1;

START1:PROCESS(CLK_100,RUN)
BEGIN
	IF(RUNIN'EVENT AND RUNIN='1') THEN
		IF(MODE_NUM="000" AND SET_NUM="110") THEN
			START<=NOT START;
		END IF;
	END IF;
END PROCESS START1;

CLR1:PROCESS(CLK_100,CLRIN)
BEGIN
	IF(CLRIN='1') THEN
		CLR<='1';
	ELSE
		CLR<='0';
	END IF;
END PROCESS CLR1;

EDIT:PROCESS(ADD,START)
BEGIN
	IF(MODE_NUM="001" AND START='0' AND CLR='0' AND SET_NUM="110") THEN
		CAL_E0R<=CAL_D0;
		CAL_E1R<=CAL_D1;
		CAL_E2R<=CAL_D2;
		CAL_E3R<=CAL_D3;
		CAL_E4R<=CAL_D4;
		CAL_E5R<=CAL_D5;
	ELSIF(MODE_NUM="001" AND CLR='1' AND START='0') THEN
		CAL_E0R<="0000";
		CAL_E1R<="0000";
		CAL_E2R<="0000";
		CAL_E3R<="0000";
		CAL_E4R<="0000";
		CAL_E5R<="0000";
	ELSIF((ADD'EVENT AND ADD='1') AND SET_NUM/="110") THEN
		IF(MODE_NUM="001" AND SET_NUM="000") THEN
			IF(CAL_E0R>="1001") THEN
				CAL_E0R<="0001";
			ELSE
				CAL_E0R<=CAL_E0R+1;
			END IF;

		ELSIF(MODE_NUM="001" AND SET_NUM="001") THEN
			IF(CAL_E1R>="0011") THEN
				CAL_E1R<="0000";
			ELSE
				CAL_E1R<=CAL_E1R+1;
			END IF;

		ELSIF(MODE_NUM="001" AND SET_NUM="010") THEN
			IF(CAL_E2R>="1001") THEN
				CAL_E2R<="0001";
			ELSE
				CAL_E2R<=CAL_E2R+1;
			END IF;

		ELSIF(MODE_NUM="001" AND SET_NUM="011") THEN
			IF(CAL_E3R>="0001") THEN
				CAL_E3R<="0000";
			ELSE
				CAL_E3R<=CAL_E3R+1;
			END IF;

		ELSIF(MODE_NUM="001" AND SET_NUM="100") THEN
			IF(CAL_E4R>="1001") THEN
				CAL_E4R<="0000";
			ELSE
				CAL_E4R<=CAL_E4R+1;
			END IF;

		ELSIF(MODE_NUM="001" AND SET_NUM="101") THEN
			IF(CAL_E5R>="1001") THEN
				CAL_E5R<="0000";
			ELSE
				CAL_E5R<=CAL_E5R+1;
			END IF;
		END IF;
	END IF;
END PROCESS EDIT;

RUN2:PROCESS(CLK_100,CAL_ADD)
BEGIN
	IF(START='1') THEN
		IF(CAL_ADD'EVENT AND CAL_ADD='1') THEN
			IF(CAL_D0R>="1001") THEN
				CAL_D0R<="0001";
				CAL_D1R<=CAL_D1R+1;
				
				IF(CAL_D1R>="0011") THEN
					CAL_D1R<="0000";
					CAL_D2R<=CAL_D2R+1;
					
					IF(CAL_D2R>="1001") THEN
						CAL_D2R<="0000";
						CAL_D3R<=CAL_D3R+1;
						
						IF(CAL_D3R>="0001") THEN
							CAL_D3R<="0000";
							CAL_D4R<=CAL_D4R+1;
							
							IF(CAL_D4R>="0010") THEN
								CAL_D4R<="0000";
								CAL_D5R<=CAL_D5R+1;
								
								IF(CAL_D5R>="1001") THEN
									CAL_D5R<="0000";
								END IF;
							END IF;
						END IF;
					END IF;
				END IF;
			ELSE
				CAL_D0R<=CAL_D0R+1;
			END IF;
		END IF;
	ELSIF(MODE_NUM="001" AND START='0') THEN
		CAL_D0R<=CAL_E0;
		CAL_D1R<=CAL_E1;
		CAL_D2R<=CAL_E2;
		CAL_D3R<=CAL_E3;
		CAL_D4R<=CAL_E4;
		CAL_D5R<=CAL_E5;
	END IF;
END PROCESS RUN2;

END ARCHITECTURE BEHAVE;