LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_UNSIGNED.ALL;

ENTITY DIV_HZ IS
PORT(
	CLK_50M: IN STD_LOGIC;		--板载晶振50MHz输入
	CLK_1: BUFFER STD_LOGIC;	--1Hz信号输出，用于秒进位
	CLK_2: BUFFER STD_LOGIC;	--2Hz信号输出，用于选定闪烁
	CLK_100: BUFFER STD_LOGIC;	--100Hz信号输出，用于百分秒进位
	CLK_800: BUFFER STD_LOGIC;	--800Hz信号输出，用于数码管动态扫描
	CLK_20K: BUFFER STD_LOGIC);	--20kHz信号输出，用于消抖按键扫描

END ENTITY DIV_HZ;

ARCHITECTURE DIV OF DIV_HZ IS
SIGNAL F1: INTEGER RANGE 0 TO 25000000;
SIGNAL F2: INTEGER RANGE 0 TO 12500000;
SIGNAL F100: INTEGER RANGE 0 TO 250000;
SIGNAL F800: INTEGER RANGE 0 TO 31250;
SIGNAL F20K: INTEGER RANGE 0 TO 1250;
	
BEGIN
DIV_1HZ:PROCESS(CLK_50M)--1Hz信号产生进程
BEGIN
	IF(CLK_50M'EVENT AND CLK_50M='1') THEN
		F1<=F1+1;
		IF (F1=25000000) THEN--当计数到2.5M时反转一次电平
			F1<=0;
			CLK_1<= NOT CLK_1;
		END IF;
	END IF;
END PROCESS DIV_1HZ;

DIV_2HZ:PROCESS(CLK_50M)--2Hz信号产生进程
BEGIN
	IF(CLK_50M'EVENT AND CLK_50M='1') THEN
		F2<=F2+1;
		IF (F2=12500000) THEN
			F2<=0;
			CLK_2<= NOT CLK_2;
		END IF;
	END IF;
END PROCESS DIV_2HZ;
	
DIV_100HZ:PROCESS(CLK_50M)--100Hz信号输出进程
BEGIN
	IF(CLK_50M'EVENT AND CLK_50M='1') THEN
		F100<=F100+1;
		IF (F100=250000) THEN
			F100<=0;
			CLK_100<= NOT CLK_100;
		END IF;
	END IF;
END PROCESS DIV_100HZ;
	
DIV_800HZ:PROCESS(CLK_50M)--800Hz信号输出进程
BEGIN
	IF(CLK_50M'EVENT AND CLK_50M='1') THEN
		F800<=F800+1;
		IF (F800=31250) THEN
			F800<=0;
			CLK_800<= NOT CLK_800;
		END IF;
	END IF;
END PROCESS DIV_800HZ;
	
DIV_20KHZ:PROCESS(CLK_50M)--20kHz信号输出进程
BEGIN
	IF(CLK_50M'EVENT AND CLK_50M='1') THEN
		F20K<=F20K+1;
		IF (F20K=1250) THEN
			F20K<=0;
			CLK_20K<= NOT CLK_20K;
		END IF;
	END IF;
END PROCESS DIV_20KHZ;

END ARCHITECTURE DIV;