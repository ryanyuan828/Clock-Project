LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_UNSIGNED.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

ENTITY ClockProject IS
PORT(
	CLK_50M:IN STD_LOGIC;--外部CLK_50K输入,用于计数产生各种频率信号输出
	BUT:IN STD_LOGIC_VECTOR(1 TO 8);--开发板按键BUT1-8
	LED:OUT STD_LOGIC_VECTOR(1 TO 8);--开发板LED灯1-8
	SEG_NCS:OUT STD_LOGIC_VECTOR(1 TO 6);--数码管选位信号
	SEG_LED:OUT STD_LOGIC_VECTOR(7 DOWNTO 0)--数码管数据信号
);
END ClockProject;

ARCHITECTURE BEHAVE OF ClockProject IS 

COMPONENT CONTROL IS
PORT(
	CLK_2,SETOUT,MODEOUT,ACKOUT: IN STD_LOGIC;--相当于按下MODE、SET等按键
	SET_NUM: INOUT STD_LOGIC_VECTOR(2 DOWNTO 0);--用于选择不同功能模块
	MODE_NUM: INOUT STD_LOGIC_VECTOR(2 DOWNTO 0);--用于选择对应位的数据
	HMS_START,STOPW_START,CAL_START,TIMER_START: IN STD_LOGIC----用于选择不同数码管信号输出
);
END COMPONENT CONTROL;

COMPONENT DEBOUNCE IS
PORT(
	CLK_2,CLK_20K: IN STD_LOGIC;--用于消抖模块扫描按键
	BUT: IN STD_LOGIC_VECTOR(1 TO 8);--用于消抖处理
	LED: OUT STD_LOGIC_VECTOR(1 TO 8);
	SETOUT,MODEOUT,CLROUT,ACKOUT,RUNOUT,ADDOUT,SUBOUT: OUT STD_LOGIC;--产生设置、模式、确认、清零、运行/暂停、加一信号
	ALM_END: IN STD_LOGIC--闹钟模块到点信号输出
);
END COMPONENT DEBOUNCE;

COMPONENT DISPLAY IS
PORT(
	CLK_1,CLK_2,CLK_800: IN STD_LOGIC;--用于数码管点闪烁、选位闪烁、动态扫描
	DIS_OUT: OUT STD_LOGIC_VECTOR(7 DOWNTO 0);--数码管数据信号
	DIS_BIT_SEL_OUT: OUT STD_LOGIC_VECTOR(5 DOWNTO 0);--数码管选位信号
	
	HMS_E5,HMS_E4,HMS_E3,HMS_E2,HMS_E1,HMS_E0: IN STD_LOGIC_VECTOR(3 DOWNTO 0);
	HMS_D5,HMS_D4,HMS_D3,HMS_D2,HMS_D1,HMS_D0: IN STD_LOGIC_VECTOR(3 DOWNTO 0);
	
	CAL_E5,CAL_E4,CAL_E3,CAL_E2,CAL_E1,CAL_E0: IN STD_LOGIC_VECTOR(3 DOWNTO 0);
	CAL_D5,CAL_D4,CAL_D3,CAL_D2,CAL_D1,CAL_D0: IN STD_LOGIC_VECTOR(3 DOWNTO 0);
	
	STOPW_D5,STOPW_D4,STOPW_D3,STOPW_D2,STOPW_D1,STOPW_D0: IN STD_LOGIC_VECTOR(3 DOWNTO 0);
	
	TIMER_E5,TIMER_E4,TIMER_E3,TIMER_E2,TIMER_E1,TIMER_E0: IN STD_LOGIC_VECTOR(3 DOWNTO 0);
	TIMER_D5,TIMER_D4,TIMER_D3,TIMER_D2,TIMER_D1,TIMER_D0: IN STD_LOGIC_VECTOR(3 DOWNTO 0);
	
	ALM_E5,ALM_E4,ALM_E3,ALM_E2,ALM_E1,ALM_E0: IN STD_LOGIC_VECTOR(3 DOWNTO 0);
	ALM_D5,ALM_D4,ALM_D3,ALM_D2,ALM_D1,ALM_D0: IN STD_LOGIC_VECTOR(3 DOWNTO 0);
	--各个模块修改、显示模式数据输出
	MODE_NUM: IN STD_LOGIC_VECTOR(2 DOWNTO 0);--用于选择不同功能模块
	SET_NUM: IN STD_LOGIC_VECTOR(2 DOWNTO 0);--用于选择对应位的数据
	HMS_START,STOPW_START,CAL_START,TIMER_START: IN STD_LOGIC;--用于选择不同数码管信号输出
	TIMER_FINISH,ALM_START: IN STD_LOGIC--用于选择对应位的数据
);
END COMPONENT DISPLAY;

COMPONENT DIV_HZ IS
PORT(
	CLK_50M: IN STD_LOGIC;--用于计数产生各种频率信号输出
	CLK_1: BUFFER STD_LOGIC;--产生1Hz信号，用于时钟模块秒进位
	CLK_2: BUFFER STD_LOGIC;--产生2Hz信号，用于数码管选位闪烁
	CLK_100: BUFFER STD_LOGIC;--产生100Hz信号，用于秒表百分位进位
	CLK_800: BUFFER STD_LOGIC;--产生800Hz信号，用于数码管动态扫描
	CLK_20K: BUFFER STD_LOGIC--产生20kHz信号，用于消抖模块扫描按键
);
END COMPONENT DIV_HZ;

COMPONENT HMS IS
PORT(
	CLK_1,CLK_100:IN STD_LOGIC;--用于时钟模块秒进位、模块内进程运行
	SETIN,CLRIN,RUNIN,ADDIN: IN STD_LOGIC;--按键消抖后信号输入
	SET_NUM:IN STD_LOGIC_VECTOR(2 DOWNTO 0);--用于选择对应位的数据块
	MODE_NUM: IN STD_LOGIC_VECTOR(2 DOWNTO 0);--用于选择不同功能模
	
	HMS_E5,HMS_E4,HMS_E3,HMS_E2,HMS_E1,HMS_E0: INOUT STD_LOGIC_VECTOR(3 DOWNTO 0);
	HMS_D5,HMS_D4,HMS_D3,HMS_D2,HMS_D1,HMS_D0: INOUT STD_LOGIC_VECTOR(3 DOWNTO 0);
	HMS_START: OUT STD_LOGIC;--时钟模式运行状态输出
	CAL_ADD:OUT STD_LOGIC--日历模式进位信号输出
);
END COMPONENT HMS;

COMPONENT CALENDAR IS
PORT(
	CLK_100:IN STD_LOGIC;--模块内进程运行
	SETIN,CLRIN,RUNIN,ADDIN: IN STD_LOGIC;--按键消抖后信号输入
	SET_NUM:IN STD_LOGIC_VECTOR(2 DOWNTO 0);--用于选择对应位的数据块
	MODE_NUM: IN STD_LOGIC_VECTOR(2 DOWNTO 0);--用于选择不同功能模式
	
	CAL_E5,CAL_E4,CAL_E3,CAL_E2,CAL_E1,CAL_E0: INOUT STD_LOGIC_VECTOR(3 DOWNTO 0);
	CAL_D5,CAL_D4,CAL_D3,CAL_D2,CAL_D1,CAL_D0: INOUT STD_LOGIC_VECTOR(3 DOWNTO 0);
	CAL_START: OUT STD_LOGIC;--日历模式运行状态输出
	CAL_ADD: IN STD_LOGIC--日历模式进位信号输入
);
END COMPONENT CALENDAR;

COMPONENT STOPWATCH IS
PORT(
	CLK_100: IN STD_LOGIC;
	RUNIN,CLRIN: IN STD_LOGIC;
	MODE_NUM: IN STD_lOGIC_VECTOR(2 DOWNTO 0);
	STOPW_D5,STOPW_D4,STOPW_D3,STOPW_D2,STOPW_D1,STOPW_D0: BUFFER STD_LOGIC_VECTOR(3 DOWNTO 0);
	STOPW_START: OUT STD_LOGIC--秒表模式运行状态输出
);
END COMPONENT STOPWATCH;

COMPONENT TIMER IS
PORT(
	CLK_1,CLK_100:IN STD_LOGIC;
	SETIN,CLRIN,RUNIN,ADDIN: IN STD_LOGIC;
	SET_NUM:IN STD_LOGIC_VECTOR(2 DOWNTO 0);
	MODE_NUM: IN STD_LOGIC_VECTOR(2 DOWNTO 0);
	
	TIMER_E5,TIMER_E4,TIMER_E3,TIMER_E2,TIMER_E1,TIMER_E0: INOUT STD_LOGIC_VECTOR(3 DOWNTO 0);
	TIMER_D5,TIMER_D4,TIMER_D3,TIMER_D2,TIMER_D1,TIMER_D0: INOUT STD_LOGIC_VECTOR(3 DOWNTO 0);
	TIMER_START,TIMER_FINISH: OUT STD_LOGIC--倒计时模式运行状态、结束状态输出
);
END COMPONENT TIMER;

COMPONENT ALARM IS
PORT(
	CLK_100:IN STD_LOGIC;
	SETIN,CLRIN,RUNIN,ADDIN: IN STD_LOGIC;
	SET_NUM:IN STD_LOGIC_VECTOR(2 DOWNTO 0);
	MODE_NUM: IN STD_LOGIC_VECTOR(2 DOWNTO 0);		--用于判断设置的闹钟时间与现在时钟模式的时间
	HMS_E5,HMS_E4,HMS_E3,HMS_E2,HMS_E1,HMS_E0: IN STD_LOGIC_VECTOR(3 DOWNTO 0);
	HMS_D5,HMS_D4,HMS_D3,HMS_D2,HMS_D1,HMS_D0: IN STD_LOGIC_VECTOR(3 DOWNTO 0);
	ALM_E5,ALM_E4,ALM_E3,ALM_E2,ALM_E1,ALM_E0: INOUT STD_LOGIC_VECTOR(3 DOWNTO 0);
	ALM_D5,ALM_D4,ALM_D3,ALM_D2,ALM_D1,ALM_D0: INOUT STD_LOGIC_VECTOR(3 DOWNTO 0);
	ALM_START,ALM_END: OUT STD_LOGIC;
	BUT6: IN STD_LOGIC
);
END COMPONENT ALARM;

SIGNAL CLK_1,CLK_2,CLK_100,CLK_800,CLK_20K: STD_LOGIC;
SIGNAL SETOUT,MODEOUT,CLROUT,ACKOUT,RUNOUT,ADDOUT,SUBOUT,BLANK: STD_LOGIC;
SIGNAL HMS_E5,HMS_E4,HMS_E3,HMS_E2,HMS_E1,HMS_E0: STD_LOGIC_VECTOR(3 DOWNTO 0);
SIGNAL HMS_D5,HMS_D4,HMS_D3,HMS_D2,HMS_D1,HMS_D0: STD_LOGIC_VECTOR(3 DOWNTO 0);

SIGNAL CAL_E5,CAL_E4,CAL_E3,CAL_E2,CAL_E1,CAL_E0: STD_LOGIC_VECTOR(3 DOWNTO 0);
SIGNAL CAL_D5,CAL_D4,CAL_D3,CAL_D2,CAL_D1,CAL_D0: STD_LOGIC_VECTOR(3 DOWNTO 0);

SIGNAL STOPW_D5,STOPW_D4,STOPW_D3,STOPW_D2,STOPW_D1,STOPW_D0: STD_LOGIC_VECTOR(3 DOWNTO 0);

SIGNAL TIMER_E5,TIMER_E4,TIMER_E3,TIMER_E2,TIMER_E1,TIMER_E0: STD_LOGIC_VECTOR(3 DOWNTO 0);
SIGNAL TIMER_D5,TIMER_D4,TIMER_D3,TIMER_D2,TIMER_D1,TIMER_D0: STD_LOGIC_VECTOR(3 DOWNTO 0);

SIGNAL ALM_E5,ALM_E4,ALM_E3,ALM_E2,ALM_E1,ALM_E0: STD_LOGIC_VECTOR(3 DOWNTO 0);
SIGNAL ALM_D5,ALM_D4,ALM_D3,ALM_D2,ALM_D1,ALM_D0: STD_LOGIC_VECTOR(3 DOWNTO 0);

SIGNAL SETIN,MODEIN,CLRIN,ACKIN,RUNIN,ADDIN,SUBIN: STD_LOGIC;
SIGNAL SET_NUM: STD_LOGIC_VECTOR(2 DOWNTO 0):="110";
SIGNAL MODE_NUM: STD_LOGIC_VECTOR(2 DOWNTO 0):="000";
SIGNAL HMS_START,CAL_START,CAL_ADD,STOPW_START,TIMER_START,TIMER_FINISH: STD_LOGIC;
SIGNAL ALM_START,ALM_END,BUT6: STD_LOGIC;

BEGIN
DIV:DIV_HZ PORT MAP(CLK_50M,CLK_1,CLK_2,CLK_100,CLK_800,CLK_20K);

DEB:DEBOUNCE PORT MAP(CLK_2,CLK_20K,BUT(1 TO 8),LED(1 TO 8),
	SETOUT,MODEOUT,CLROUT,ACKOUT,RUNOUT,ADDOUT,SUBOUT,ALM_END);

CON:CONTROL PORT MAP(
	CLK_2,SETOUT,MODEOUT,ACKOUT,SET_NUM,MODE_NUM,
	HMS_START,STOPW_START,CAL_START,TIMER_START);
	
DIS:DISPLAY PORT MAP(
	CLK_1,CLK_2,CLK_800,SEG_LED(7 DOWNTO 0),SEG_NCS(1 TO 6),
	HMS_E5,HMS_E4,HMS_E3,HMS_E2,HMS_E1,HMS_E0,
	HMS_D5,HMS_D4,HMS_D3,HMS_D2,HMS_D1,HMS_D0,
	CAL_E5,CAL_E4,CAL_E3,CAL_E2,CAL_E1,CAL_E0,
	CAL_D5,CAL_D4,CAL_D3,CAL_D2,CAL_D1,CAL_D0,
	STOPW_D5,STOPW_D4,STOPW_D3,STOPW_D2,STOPW_D1,STOPW_D0,
	TIMER_E5,TIMER_E4,TIMER_E3,TIMER_E2,TIMER_E1,TIMER_E0,
	TIMER_D5,TIMER_D4,TIMER_D3,TIMER_D2,TIMER_D1,TIMER_D0,
	ALM_E5,ALM_E4,ALM_E3,ALM_E2,ALM_E1,ALM_E0,
	ALM_D5,ALM_D4,ALM_D3,ALM_D2,ALM_D1,ALM_D0,
	MODE_NUM,SET_NUM,HMS_START,STOPW_START,CAL_START,TIMER_START,TIMER_FINISH,ALM_START);
	
SFM:HMS PORT MAP(
	CLK_1,CLK_100,SETOUT,CLROUT,RUNOUT,ADDOUT,SET_NUM,MODE_NUM,
	HMS_E5,HMS_E4,HMS_E3,HMS_E2,HMS_E1,HMS_E0,
	HMS_D5,HMS_D4,HMS_D3,HMS_D2,HMS_D1,HMS_D0,HMS_START,CAL_ADD);

CAL:CALENDAR PORT MAP(
	CLK_100,SETOUT,CLROUT,RUNOUT,ADDOUT,SET_NUM,MODE_NUM,
	CAL_E5,CAL_E4,CAL_E3,CAL_E2,CAL_E1,CAL_E0,
	CAL_D5,CAL_D4,CAL_D3,CAL_D2,CAL_D1,CAL_D0,
	CAL_START,CAL_ADD);	
	
STO:STOPWATCH PORT MAP(
	CLK_100,RUNOUT,CLROUT,MODE_NUM,STOPW_D5,STOPW_D4,STOPW_D3,STOPW_D2,STOPW_D1,STOPW_D0,STOPW_START);
	
TIM:TIMER PORT MAP(
    CLK_1,CLK_100,SETOUT,CLROUT,RUNOUT,ADDOUT,SET_NUM,MODE_NUM,
	TIMER_E5,TIMER_E4,TIMER_E3,TIMER_E2,TIMER_E1,TIMER_E0,
	TIMER_D5,TIMER_D4,TIMER_D3,TIMER_D2,TIMER_D1,TIMER_D0,TIMER_START,TIMER_FINISH);
	
ALM:ALARM PORT MAP(
	CLK_100,SETOUT,CLROUT,RUNOUT,ADDOUT,SET_NUM,MODE_NUM,
	HMS_E5,HMS_E4,HMS_E3,HMS_E2,HMS_E1,HMS_E0,
	HMS_D5,HMS_D4,HMS_D3,HMS_D2,HMS_D1,HMS_D0,
	ALM_E5,ALM_E4,ALM_E3,ALM_E2,ALM_E1,ALM_E0,
	ALM_D5,ALM_D4,ALM_D3,ALM_D2,ALM_D1,ALM_D0,
	ALM_START,ALM_END,BUT(6)
);
	
END ARCHITECTURE BEHAVE;