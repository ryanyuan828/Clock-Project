LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_UNSIGNED.ALL;

ENTITY TIMER IS
PORT(
	CLK_1,CLK_100:IN STD_LOGIC;
	SETIN,CLRIN,RUNIN,ADDIN: IN STD_LOGIC;
	SET_NUM:IN STD_LOGIC_VECTOR(2 DOWNTO 0);
	MODE_NUM: IN STD_LOGIC_VECTOR(2 DOWNTO 0);
	
	TIMER_E5,TIMER_E4,TIMER_E3,TIMER_E2,TIMER_E1,TIMER_E0: INOUT STD_LOGIC_VECTOR(3 DOWNTO 0);
	TIMER_D5,TIMER_D4,TIMER_D3,TIMER_D2,TIMER_D1,TIMER_D0: INOUT STD_LOGIC_VECTOR(3 DOWNTO 0);
	TIMER_START,TIMER_FINISH: OUT STD_LOGIC
);
END ENTITY TIMER;

ARCHITECTURE BEHAVE OF TIMER IS
SIGNAL TIMER_E5R,TIMER_E4R,TIMER_E3R,TIMER_E2R,TIMER_E1R,TIMER_E0R: STD_LOGIC_VECTOR(3 DOWNTO 0);
SIGNAL TIMER_D5R,TIMER_D4R,TIMER_D3R,TIMER_D2R,TIMER_D1R,TIMER_D0R: STD_LOGIC_VECTOR(3 DOWNTO 0);
SIGNAL START,FINISH: STD_LOGIC:='0';
SIGNAL CLR: STD_LOGIC:='1';
SIGNAL RUN,ADD: STD_LOGIC;

BEGIN
TIMER_E5<=TIMER_E5R;--将寄存的修改状态信号输出数码管
TIMER_E4<=TIMER_E4R;
TIMER_E3<=TIMER_E3R;
TIMER_E2<=TIMER_E2R;
TIMER_E1<=TIMER_E1R;
TIMER_E0<=TIMER_E0R;

TIMER_D5<=TIMER_D5R;--将寄存的显示状态信号输出数码管
TIMER_D4<=TIMER_D4R;
TIMER_D3<=TIMER_D3R;
TIMER_D2<=TIMER_D2R;
TIMER_D1<=TIMER_D1R;
TIMER_D0<=TIMER_D0R;

TIMER_START<=START;
TIMER_FINISH<=FINISH;

ADD1:PROCESS(ADDIN)
BEGIN
	IF(MODE_NUM="011" AND ADDIN='1') THEN
		ADD<='1';--在倒计时模式下按ADD键才可以加一
	ELSE
		ADD<='0';
	END IF;
END PROCESS ADD1;

START1:PROCESS(CLK_100,RUNIN)
BEGIN
	IF(MODE_NUM="011" AND SET_NUM="110") THEN
		IF(RUNIN'EVENT AND RUNIN='1') THEN
			START<=NOT START;--在倒计时模式下按RUN键切换运行状态
		END IF;
		
		IF(START='1' AND (TIMER_D5="0000" AND TIMER_D4="0000" AND TIMER_D3="0000" AND TIMER_D2="0000" AND TIMER_D1="0000" AND TIMER_D0="0000")) THEN
			FINISH<='1';--当所有显示状态的数码管数据为0时输出结束信号
		ELSE
			FINISH<='0';
		END IF;
	END IF;
END PROCESS START1;

CLR1:PROCESS(CLRIN)
BEGIN
	IF(CLRIN='1') THEN
		CLR<='1';--当按下CLR键清零
	ELSE
		CLR<='0';
	END IF;
END PROCESS CLR1;

EDIT:PROCESS(ADD,START)--手动修改模式
BEGIN
	IF(MODE_NUM="011" AND START='0' AND CLR='0' AND SET_NUM="110") THEN
		TIMER_E0R<=TIMER_D0;
		TIMER_E1R<=TIMER_D1;
		TIMER_E2R<=TIMER_D2;
		TIMER_E3R<=TIMER_D3;
		TIMER_E4R<=TIMER_D4;
		TIMER_E5R<=TIMER_D5;
	ELSIF(MODE_NUM="011" AND CLR='1') THEN
		TIMER_E0R<="0000";
		TIMER_E1R<="0000";
		TIMER_E2R<="0000";
		TIMER_E3R<="0000";
		TIMER_E4R<="0000";
		TIMER_E5R<="0000";
	ELSIF((ADD'EVENT AND ADD='1') AND SET_NUM/="110") THEN
		IF(MODE_NUM="011" AND SET_NUM="000") THEN
			IF(TIMER_E0R>="1001") THEN
				TIMER_E0R<="0000";
			ELSE
				TIMER_E0R<=TIMER_E0R+1;
			END IF;

		ELSIF(MODE_NUM="011" AND SET_NUM="001") THEN
			IF(TIMER_E1R>="0101") THEN
				TIMER_E1R<="0000";
			ELSE
				TIMER_E1R<=TIMER_E1R+1;
			END IF;

		ELSIF(MODE_NUM="011" AND SET_NUM="010") THEN
			IF(TIMER_E2R>="1001") THEN
				TIMER_E2R<="0000";
			ELSE
				TIMER_E2R<=TIMER_E2R+1;
			END IF;

		ELSIF(MODE_NUM="011" AND SET_NUM="011") THEN
			IF(TIMER_E3R>="0101") THEN
				TIMER_E3R<="0000";
			ELSE
				TIMER_E3R<=TIMER_E3R+1;
			END IF;

		ELSIF(MODE_NUM="011" AND SET_NUM="100") THEN
			IF(TIMER_E4R>="1001") THEN
				TIMER_E4R<="0000";
			ELSE
				TIMER_E4R<=TIMER_E4R+1;
			END IF;

		ELSIF(MODE_NUM="011" AND SET_NUM="101") THEN
			IF(TIMER_E5R>="1001") THEN
				TIMER_E5R<="0000";
			ELSE
				TIMER_E5R<=TIMER_E5R+1;
			END IF;
		END IF;
	END IF;
END PROCESS EDIT;

RUN2:PROCESS(CLK_100,CLK_1)
BEGIN
	IF(CLK_1'EVENT AND CLK_1='1') THEN
		IF(START='1' AND FINISH='0') THEN
			IF(TIMER_D0R="0000") THEN
				TIMER_D0R<="1001";
				TIMER_D1R<=TIMER_D1R-1;
				
				IF(TIMER_D1R="0000") THEN
					TIMER_D1R<="0101";
					TIMER_D2R<=TIMER_D2R-1;
					
					IF(TIMER_D2R="0000") THEN
						TIMER_D2R<="1001";
						TIMER_D3R<=TIMER_D3R-1;
						
						IF(TIMER_D3R="0000") THEN
							TIMER_D3R<="0101";
							TIMER_D4R<=TIMER_D4R-1;
							
							IF(TIMER_D4R="0000") THEN
								TIMER_D4R<="1001";
								TIMER_D5R<=TIMER_D5R-1;
							END IF;
						END IF;
					END IF;
				END IF;
			ELSE
				TIMER_D0R<=TIMER_D0R-1;
			END IF;
		ELSIF(MODE_NUM="011" AND START='0') THEN
			TIMER_D0R<=TIMER_E0;
			TIMER_D1R<=TIMER_E1;
			TIMER_D2R<=TIMER_E2;
			TIMER_D3R<=TIMER_E3;
			TIMER_D4R<=TIMER_E4;
			TIMER_D5R<=TIMER_E5;
		END IF;
	END IF;
END PROCESS RUN2;

END ARCHITECTURE BEHAVE;