LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_UNSIGNED.ALL;

ENTITY HMS IS
PORT(
	CLK_1,CLK_100:IN STD_LOGIC;
	SETIN,CLRIN,RUNIN,ADDIN: IN STD_LOGIC;
	SET_NUM:IN STD_LOGIC_VECTOR(2 DOWNTO 0);
	MODE_NUM: IN STD_LOGIC_VECTOR(2 DOWNTO 0);
	
	HMS_E5,HMS_E4,HMS_E3,HMS_E2,HMS_E1,HMS_E0: INOUT STD_LOGIC_VECTOR(3 DOWNTO 0);
	HMS_D5,HMS_D4,HMS_D3,HMS_D2,HMS_D1,HMS_D0: INOUT STD_LOGIC_VECTOR(3 DOWNTO 0);
	HMS_START: OUT STD_LOGIC;--输出运行状态
	CAL_ADD:OUT STD_LOGIC--日历模块进位信号输出，实现与日历模块联动
);
END ENTITY HMS;

ARCHITECTURE BEHAVE OF HMS IS
SIGNAL HMS_E5R,HMS_E4R,HMS_E3R,HMS_E2R,HMS_E1R,HMS_E0R: STD_LOGIC_VECTOR(3 DOWNTO 0);
SIGNAL HMS_D5R,HMS_D4R,HMS_D3R,HMS_D2R,HMS_D1R,HMS_D0R: STD_LOGIC_VECTOR(3 DOWNTO 0);
SIGNAL START: STD_LOGIC:='0';
SIGNAL CLR: STD_LOGIC:='1';
SIGNAL RUN,ADD: STD_LOGIC;

BEGIN
HMS_E5<=HMS_E5R;--将寄存的修改状态信号输出数码管
HMS_E4<=HMS_E4R;
HMS_E3<=HMS_E3R;
HMS_E2<=HMS_E2R;
HMS_E1<=HMS_E1R;
HMS_E0<=HMS_E0R;

HMS_D5<=HMS_D5R;--将寄存的显示状态信号输出数码管
HMS_D4<=HMS_D4R;
HMS_D3<=HMS_D3R;
HMS_D2<=HMS_D2R;
HMS_D1<=HMS_D1R;
HMS_D0<=HMS_D0R;
HMS_START<=START;

ADD1:PROCESS(ADDIN)
BEGIN
	IF(MODE_NUM="000" AND ADDIN='1') THEN
		ADD<='1';--在时钟模式下按ADD键才可以加一
	ELSE
		ADD<='0';
	END IF;
END PROCESS ADD1;

START1:PROCESS(CLK_100,RUN)
BEGIN
	IF(RUNIN'EVENT AND RUNIN='1') THEN
		IF(MODE_NUM="000" AND SET_NUM="110") THEN
			START<=NOT START;--在时钟模式下按RUN键切换运行状态
		END IF;
	END IF;
END PROCESS START1;

CLR1:PROCESS(CLRIN)
BEGIN
	IF(CLRIN='1') THEN
		CLR<='1';--当按下CLR键清零
	ELSE
		CLR<='0';
	END IF;
END PROCESS CLR1;

EDIT:PROCESS(ADD,START)--手动修改模式
BEGIN--当在时钟模式且不在运行状态且没有按下CLR键，将显示状态数据传给修改状态寄存
	IF(MODE_NUM="000" AND START='0' AND CLR='0' AND SET_NUM="110") THEN
		HMS_E0R<=HMS_D0;
		HMS_E1R<=HMS_D1;
		HMS_E2R<=HMS_D2;
		HMS_E3R<=HMS_D3;
		HMS_E4R<=HMS_D4;
		HMS_E5R<=HMS_D5;
	ELSIF(MODE_NUM="000" AND CLR='1' AND START='0') THEN
		HMS_E0R<="0000";--当在时钟模式且按下CLR键且不在运行状态时才可清零
		HMS_E1R<="0000";
		HMS_E2R<="0000";
		HMS_E3R<="0000";
		HMS_E4R<="0000";
		HMS_E5R<="0000";--当在时钟模式且按下ADD键，给对应数码管加一
	ELSIF((ADD'EVENT AND ADD='1') AND SET_NUM/="110") THEN
		IF(MODE_NUM="000" AND SET_NUM="000") THEN
			IF(HMS_E0R>="1001") THEN
				HMS_E0R<="0000";--当加一后超过9设为0
			ELSE
				HMS_E0R<=HMS_E0R+1;
			END IF;

		ELSIF(MODE_NUM="000" AND SET_NUM="001") THEN
			IF(HMS_E1R>="0101") THEN
				HMS_E1R<="0000";--当加一后超过6设为0
			ELSE
				HMS_E1R<=HMS_E1R+1;
			END IF;

		ELSIF(MODE_NUM="000" AND SET_NUM="010") THEN
			IF(HMS_E2R>="1001") THEN
				HMS_E2R<="0000";--当加一后超过9设为0
			ELSE
				HMS_E2R<=HMS_E2R+1;
			END IF;

		ELSIF(MODE_NUM="000" AND SET_NUM="011") THEN
			IF(HMS_E3R>="0101") THEN
				HMS_E3R<="0000";--当加一后超过6设为0
			ELSE
				HMS_E3R<=HMS_E3R+1;
			END IF;

		ELSIF(MODE_NUM="000" AND SET_NUM="100") THEN
			IF(HMS_E4R>="1001") THEN
				HMS_E4R<="0000";--当加一后超过9设为0
			ELSE
				HMS_E4R<=HMS_E4R+1;
			END IF;

		ELSIF(MODE_NUM="000" AND SET_NUM="101") THEN
			IF(HMS_E5R>="0010") THEN
				HMS_E5R<="0000";--当加一后超过2设为0
			ELSE
				HMS_E5R<=HMS_E5R+1;
			END IF;
		END IF;
	END IF;
END PROCESS EDIT;

RUN2:PROCESS(CLK_100,CLK_1)--自动运行状态
BEGIN
	IF(CLK_1'EVENT AND CLK_1='1') THEN--按1Hz频率自动加一和进位
		IF(START='1') THEN
			IF(HMS_D0R>="1001") THEN--当秒低位超过9后设为0
				HMS_D0R<="0000";
				HMS_D1R<=HMS_D1R+1;--秒高位进位
				
				IF(HMS_D1R>="0101") THEN--当秒高位超过5后设为0
					HMS_D1R<="0000";
					HMS_D2R<=HMS_D2R+1;--分低位进位
					
					IF(HMS_D2R>="1001") THEN--当分低位超过9后设为0
						HMS_D2R<="0000";
						HMS_D3R<=HMS_D3R+1;--分高位进位
						
						IF(HMS_D3R>="0101") THEN--当分高位超过5后设为0
							HMS_D3R<="0000";
							
							IF(HMS_D5R>="0010" AND HMS_D4R="0011") THEN
								HMS_D5R<="0000";--当时超过23后设为00
								HMS_D4R<="0000";
								
								CAL_ADD<='1';--同时给日历模块进位信号
								
							ELSIF(HMS_D4R>="1001") THEN--当时高位不为2且时地位超过9
								HMS_D4R<="0000";--时低位设为0
								HMS_D5R<=HMS_D5R+1;--时高位进位
							ELSE
								HMS_D4R<=HMS_D4R+1;--否则时低位进位
							END IF;
						END IF;
					END IF;
				END IF;
			ELSE
				HMS_D0R<=HMS_D0R+1;--秒低位进位
				CAL_ADD<='0';--取消日历进位信号
				
			END IF;
		ELSIF(MODE_NUM="000" AND START='0') THEN--当在时钟模式且不在运行状态
			HMS_D0R<=HMS_E0;--将修改状态的数据传给显示状态寄存器
			HMS_D1R<=HMS_E1;
			HMS_D2R<=HMS_E2;
			HMS_D3R<=HMS_E3;
			HMS_D4R<=HMS_E4;
			HMS_D5R<=HMS_E5;
		END IF;
	END IF;
END PROCESS RUN2;

END ARCHITECTURE BEHAVE;