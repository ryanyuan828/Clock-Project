LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_UNSIGNED.ALL;

ENTITY DEBOUNCE IS
PORT(
	CLK_2,CLK_20K: IN STD_LOGIC;
	BUT: IN STD_LOGIC_VECTOR(1 TO 8);
	LED: OUT STD_LOGIC_VECTOR(1 TO 8);
	SETOUT,MODEOUT,CLROUT,ACKOUT,RUNOUT,ADDOUT,SUBOUT: OUT STD_LOGIC;
	ALM_END: IN STD_LOGIC
);
END ENTITY DEBOUNCE;

ARCHITECTURE BEHAVE OF DEBOUNCE IS
SIGNAL COUNT1: INTEGER RANGE 0 TO 200:=0;
SIGNAL COUNT2: INTEGER RANGE 0 TO 200:=0;
SIGNAL COUNT3: INTEGER RANGE 0 TO 200:=0;
SIGNAL COUNT4: INTEGER RANGE 0 TO 200:=0;
SIGNAL COUNT5: INTEGER RANGE 0 TO 200:=0;
SIGNAL COUNT7: INTEGER RANGE 0 TO 200:=0;
SIGNAL COUNT8: INTEGER RANGE 0 TO 200:=0;

BEGIN
SET:PROCESS(CLK_20K,BUT)
BEGIN
	IF(BUT="01111111") THEN--当按下第1个按键
		IF(CLK_20K'EVENT AND CLK_20K='1') THEN
			IF(COUNT1=200) THEN
				COUNT1<=COUNT1;
			ELSE
				COUNT1<=COUNT1+1;
			END IF;
			
			IF(COUNT1=199) THEN--累计计数到199次（约1ms）
				SETOUT<='1';
				
			ELSE
				SETOUT<='0';--输出SETOUT高电平
				
			END IF;
		END IF;
		LED(1)<='0';
	ELSE
		COUNT1<=0;
		SETOUT<='0';
		LED(1)<='1';
	END IF;
END PROCESS SET;
	
MODE:PROCESS(CLK_20K,BUT)
BEGIN
	IF(BUT="10111111") THEN--当按下第2个按键
		IF(CLK_20K'EVENT AND CLK_20K='1') THEN
			IF(COUNT2=200) THEN
				COUNT2<=COUNT2;
			ELSE
				COUNT2<=COUNT2+1;
			END IF;
			
			IF(COUNT2=199) THEN
				MODEOUT<='1';
			ELSE
				MODEOUT<='0';
			END IF;
		END IF;
		LED(2)<='0';
	ELSE
		COUNT2<=0;
		MODEOUT<='0';
		LED(2)<='1';
	END IF;
END PROCESS MODE;

ACK:PROCESS(CLK_20K,BUT)
BEGIN
	IF(BUT="11011111") THEN--当按下第3个按键
		IF(CLK_20K'EVENT AND CLK_20K='1') THEN
			IF(COUNT3=200) THEN
				COUNT3<=COUNT3;
			ELSE
				COUNT3<=COUNT3+1;
			END IF;
			
			IF(COUNT3=199) THEN
				ACKOUT<='1';
			ELSE
				ACKOUT<='0';
			END IF;
		END IF;
		LED(3)<='0';
	ELSE
		COUNT3<=0;
		ACKOUT<='0';
		LED(3)<='1';
	END IF;
END PROCESS ACK;

CLR:PROCESS(CLK_20K,BUT)
BEGIN
	IF(BUT="11101111") THEN--当按下第4个按键
		IF(CLK_20K'EVENT AND CLK_20K='1') THEN
			IF(COUNT4=200) THEN
				COUNT4<=COUNT4;
			ELSE
				COUNT4<=COUNT4+1;
			END IF;
			
			IF(COUNT4=199) THEN
				CLROUT<='1';
			ELSE
				CLROUT<='0';
			END IF;
		END IF;
		LED(4)<='0';
	ELSE
		COUNT4<=0;
		CLROUT<='0';
		LED(4)<='1';
	END IF;
END PROCESS CLR;
	
RUN:PROCESS(CLK_20K,BUT)
BEGIN
	IF(BUT="11110111") THEN--当按下第5个按键
		IF(CLK_20K'EVENT AND CLK_20K='1') THEN
			IF(COUNT5=200) THEN
				COUNT5<=COUNT5;
			ELSE
				COUNT5<=COUNT5+1;
			END IF;
			
			IF(COUNT5=199) THEN
				RUNOUT<='1';
			ELSE
				RUNOUT<='0';
			END IF;
		END IF;
		LED(5)<='0';
	ELSE
		COUNT5<=0;
		RUNOUT<='0';
		LED(5)<='1';
	END IF;
END PROCESS RUN;

ALARM:PROCESS(CLK_2)
BEGIN
	IF(CLK_2='1') THEN--当闹钟到点时闪灯
		IF(ALM_END='1') THEN
			LED(6)<='0';
		ELSE
			LED(6)<='1';
		END IF;
	ELSE
		LED(6)<='1';
	END IF;
END PROCESS ALARM;

ADD:PROCESS(CLK_20K,BUT)
BEGIN
	IF(BUT="11111101") THEN--当按下第7个按键
		IF(CLK_20K'EVENT AND CLK_20K='1') THEN
			IF(COUNT7=200) THEN
				COUNT7<=COUNT7;
			ELSE
				COUNT7<=COUNT7+1;
			END IF;
			
			IF(COUNT7=199) THEN
				ADDOUT<='1';
			ELSE
				ADDOUT<='0';
			END IF;
		END IF;
		LED(7)<='0';
	ELSE
		COUNT7<=0;
		ADDOUT<='0';
		LED(7)<='1';
	END IF;
END PROCESS ADD;
	
SUB:PROCESS(CLK_20K,BUT)
BEGIN
	IF(BUT="11111110") THEN--当按下第8个按键
		IF(CLK_20K'EVENT AND CLK_20K='1') THEN
			IF(COUNT8=200) THEN
				COUNT8<=COUNT8;
			ELSE
				COUNT8<=COUNT8+1;
			END IF;
			
			IF(COUNT8=199) THEN
				SUBOUT<='1';
			ELSE
				SUBOUT<='0';
			END IF;
		END IF;
		LED(8)<='0';
	ELSE
		COUNT8<=0;
		SUBOUT<='0';
		LED(8)<='1';
	END IF;
END PROCESS SUB;

END ARCHITECTURE BEHAVE;