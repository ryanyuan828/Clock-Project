LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_UNSIGNED.ALL;

ENTITY ALARM IS
PORT(
	CLK_100:IN STD_LOGIC;
	SETIN,CLRIN,RUNIN,ADDIN: IN STD_LOGIC;
	SET_NUM:IN STD_LOGIC_VECTOR(2 DOWNTO 0);
	MODE_NUM: IN STD_LOGIC_VECTOR(2 DOWNTO 0);
	HMS_E5,HMS_E4,HMS_E3,HMS_E2,HMS_E1,HMS_E0: IN STD_LOGIC_VECTOR(3 DOWNTO 0);--获得时间模块当前时间
	HMS_D5,HMS_D4,HMS_D3,HMS_D2,HMS_D1,HMS_D0: IN STD_LOGIC_VECTOR(3 DOWNTO 0);
	ALM_E5,ALM_E4,ALM_E3,ALM_E2,ALM_E1,ALM_E0: INOUT STD_LOGIC_VECTOR(3 DOWNTO 0);
	ALM_D5,ALM_D4,ALM_D3,ALM_D2,ALM_D1,ALM_D0: INOUT STD_LOGIC_VECTOR(3 DOWNTO 0);
	ALM_START,ALM_END: OUT STD_LOGIC;
	BUT6: IN STD_LOGIC
);
END ENTITY ALARM;

ARCHITECTURE BEHAVE OF ALARM IS
SIGNAL ALM_E5R,ALM_E4R,ALM_E3R,ALM_E2R,ALM_E1R,ALM_E0R: STD_LOGIC_VECTOR(3 DOWNTO 0);
SIGNAL ALM_D5R,ALM_D4R,ALM_D3R,ALM_D2R,ALM_D1R,ALM_D0R: STD_LOGIC_VECTOR(3 DOWNTO 0);
SIGNAL CLR: STD_LOGIC:='1';
SIGNAL RUN,ADD: STD_LOGIC;
SIGNAL START: STD_LOGIC:='0';

BEGIN
ALM_E5<=ALM_E5R;--将寄存的修改状态信号输出数码管
ALM_E4<=ALM_E4R;
ALM_E3<=ALM_E3R;
ALM_E2<=ALM_E2R;
ALM_E1<=ALM_E1R;
ALM_E0<=ALM_E0R;

ALM_D5<=ALM_D5R;--将寄存的显示状态信号输出数码管
ALM_D4<=ALM_D4R;
ALM_D3<=ALM_D3R;
ALM_D2<=ALM_D2R;
ALM_D1<=ALM_D1R;
ALM_D0<=ALM_D0R;
ALM_START<=START;

ADD1:PROCESS(ADDIN)
BEGIN
	IF(MODE_NUM="100" AND ADDIN='1') THEN
		ADD<='1';--在闹钟模式下按ADD键才可以加一
	ELSE
		ADD<='0';
	END IF;
END PROCESS ADD1;

START1:PROCESS(CLK_100,RUN)
BEGIN
	IF(RUNIN'EVENT AND RUNIN='1') THEN
		IF(MODE_NUM="100" AND SET_NUM="110") THEN
			START<=NOT START;--在闹钟模式下按RUN键切换运行状态
		END IF;
	END IF;
END PROCESS START1;

CLR1:PROCESS(CLK_100,CLRIN)
BEGIN
	IF(CLRIN='1') THEN
		CLR<='1';--当按下CLR键清零
	ELSE
		CLR<='0';
	END IF;
END PROCESS CLR1;

EDIT:PROCESS(ADD)--手动修改模式
BEGIN
	IF(MODE_NUM="100" AND START='0' AND CLR='0' AND SET_NUM="110") THEN
		ALM_E0R<=ALM_D0;
		ALM_E1R<=ALM_D1;
		ALM_E2R<=ALM_D2;
		ALM_E3R<=ALM_D3;
		ALM_E4R<=ALM_D4;
		ALM_E5R<=ALM_D5;
	ELSIF(MODE_NUM="100" AND START='0' AND CLR='1') THEN
		ALM_E0R<="0000";
		ALM_E1R<="0000";
		ALM_E2R<="0000";
		ALM_E3R<="0000";
		ALM_E4R<="0000";
		ALM_E5R<="0000";
	ELSIF((ADD'EVENT AND ADD='1') AND SET_NUM/="110") THEN
		IF(MODE_NUM="100" AND SET_NUM="000") THEN
			IF(ALM_E0R>="1001") THEN
				ALM_E0R<="0000";
			ELSE
				ALM_E0R<=ALM_E0R+1;
			END IF;

		ELSIF(MODE_NUM="100" AND SET_NUM="001") THEN
			IF(ALM_E1R>="0101") THEN
				ALM_E1R<="0000";
			ELSE
				ALM_E1R<=ALM_E1R+1;
			END IF;

		ELSIF(MODE_NUM="100" AND SET_NUM="010") THEN
			IF(ALM_E2R>="1001") THEN
				ALM_E2R<="0000";
			ELSE
				ALM_E2R<=ALM_E2R+1;
			END IF;

		ELSIF(MODE_NUM="100" AND SET_NUM="011") THEN
			IF(ALM_E3R>="0101") THEN
				ALM_E3R<="0000";
			ELSE
				ALM_E3R<=ALM_E3R+1;
			END IF;

		ELSIF(MODE_NUM="100" AND SET_NUM="100") THEN
			IF(ALM_E4R>="1001") THEN
				ALM_E4R<="0000";
			ELSE
				ALM_E4R<=ALM_E4R+1;
			END IF;

		ELSIF(MODE_NUM="100" AND SET_NUM="101") THEN
			IF(ALM_E5R>="0010") THEN
				ALM_E5R<="0000";
			ELSE
				ALM_E5R<=ALM_E5R+1;
			END IF;
		END IF;
	END IF;
END PROCESS EDIT;

RUN1:PROCESS(CLK_100)
BEGIN
	IF(MODE_NUM="100" AND START='0') THEN
		ALM_D0R<=ALM_E0;
		ALM_D1R<=ALM_E1;
		ALM_D2R<=ALM_E2;
		ALM_D3R<=ALM_E3;
		ALM_D4R<=ALM_E4;
		ALM_D5R<=ALM_E5;
	END IF;
END PROCESS RUN1;

RUN2:PROCESS(CLK_100,BUT6)
BEGIN
	IF(HMS_D0=ALM_D0 AND HMS_D1=ALM_D1 AND HMS_D2=ALM_D2 AND HMS_D3=ALM_D3 AND HMS_D4=ALM_D4 AND HMS_D5=ALM_D5) THEN
		ALM_END<='1';--与闹钟模块时间相比，相等则输出信号
	ELSIF(BUT6='0') THEN--按下BUT6后解除信号
		ALM_END<='0';
	END IF;
END PROCESS RUN2;

END ARCHITECTURE BEHAVE;