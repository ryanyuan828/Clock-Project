LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_UNSIGNED.ALL;

ENTITY CONTROL IS
PORT(
	CLK_2,SETOUT,MODEOUT,ACKOUT: IN STD_LOGIC;
	SET_NUM:INOUT STD_LOGIC_VECTOR(2 DOWNTO 0);
	MODE_NUM:INOUT STD_LOGIC_VECTOR(2 DOWNTO 0);
	HMS_START,STOPW_START,CAL_START,TIMER_START: IN STD_LOGIC
);
END ENTITY CONTROL;

ARCHITECTURE BEHAVE OF CONTROL IS
BEGIN
SET_CALC:PROCESS(CLK_2)
BEGIN
	IF(SETOUT'EVENT AND SETOUT='1') THEN
		IF(MODE_NUM="000" AND HMS_START='0') THEN--模式为时钟且不在运行时
			IF(SET_NUM>="110") THEN--可设置位选从000->110
				SET_NUM<="000";
			ELSE
				SET_NUM<=SET_NUM+1;
			END IF;
		ELSIF(MODE_NUM="001" AND CAL_START='0') THEN--模式为日历且不在运行时
			IF(SET_NUM>="110") THEN
				SET_NUM<="000";
			ELSE
				SET_NUM<=SET_NUM+1;
			END IF;
		ELSIF(MODE_NUM="011" AND TIMER_START='0') THEN--模式为倒计时且不在运行时
			IF(SET_NUM>="110") THEN
				SET_NUM<="000";
			ELSE
				SET_NUM<=SET_NUM+1;
			END IF;
		ELSIF(MODE_NUM="100") THEN--模式为闹钟且不在运行时
			IF(SET_NUM>="110") THEN
				SET_NUM<="000";
			ELSE
				SET_NUM<=SET_NUM+1;
			END IF;
		END IF;
	END IF;
	
	IF(ACKOUT='1') THEN--按下ACK键后退出设置模式
		SET_NUM<="110";
	END IF;
END PROCESS SET_CALC;

MODE_CALC:
	PROCESS(MODEOUT)
	BEGIN
		IF(MODEOUT'EVENT AND MODEOUT='1') THEN--每按一次MODE键切换模式
			IF(MODE_NUM>="100") THEN
				MODE_NUM<="000";
			ELSE
				MODE_NUM<=MODE_NUM+1;
			END IF;
		END IF;
	END PROCESS MODE_CALC;
	
END ARCHITECTURE BEHAVE;